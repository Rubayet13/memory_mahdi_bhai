package agent_pkg;

  `include "../tb/params.sv"
  `include "mem_trans.sv"
  `include "mem_driver.sv"
  `include "mem_driver_v2.sv"
  `include "mem_monitor.sv"
  `include "mem_agent.sv"

endpackage