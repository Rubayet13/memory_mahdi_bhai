package env_pkg;

  import agent_pkg::*;
  
  `include "../tb/params.sv"
  `include "mem_scoreboard.sv"
  `include "mem_scoreboard_v2.sv"
  `include "mem_environment.sv"

endpackage