package seq_pkg;

  import agent_pkg::mem_trans;
  
  `include "../tb/params.sv"
  `include "base_seq.sv"
  `include "random_seq.sv"
  `include "write_read_seq.sv"

endpackage